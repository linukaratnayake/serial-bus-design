module split_target_port(
    input logic clk,
    input logic rst_n,
    input logic split_req,
    input logic arbiter_grant,
    input logic [7:0] target_data_out,
    input logic target_data_out_valid,
    input logic target_rw, // 1 for write, 0 for read
    input logic target_ready,
    input logic target_split_ack,
    input logic target_ack,
    input logic bus_data_in_valid,
    input logic bus_data_in,
    output logic bus_data_out,
    output logic split_grant,
    output logic [7:0] target_data_in,
    output logic target_data_in_valid,
    output logic bus_data_out_valid,
    output logic arbiter_split_req,
    output logic split_ack,
    output logic bus_target_ready,
    output logic bus_target_rw,
    output logic bus_split_ack,
    output logic bus_target_ack
);

assign split_grant = arbiter_grant;
assign arbiter_split_req = split_req;
assign bus_target_rw = target_rw;
assign bus_target_ready = target_ready;
assign bus_target_ack = target_ack;
assign bus_split_ack = target_split_ack;

logic [7:0] tx_shift;
logic [3:0] tx_bits_remaining;
logic tx_active;
logic [7:0] rx_shift;
logic [2:0] rx_bit_count;

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        tx_shift <= '0;
        tx_bits_remaining <= '0;
        tx_active <= 1'b0;
        bus_data_out <= 1'b0;
        bus_data_out_valid <= 1'b0;
    end else begin
        bus_data_out_valid <= 1'b0;

        if (tx_active) begin
            bus_data_out <= tx_shift[0];
            bus_data_out_valid <= 1'b1;
            tx_shift <= {1'b0, tx_shift[7:1]};

            if (tx_bits_remaining == 4'd1) begin
                tx_active <= 1'b0;
                tx_bits_remaining <= '0;
            end else begin
                tx_bits_remaining <= tx_bits_remaining - 4'd1;
            end
        end else if (target_data_out_valid) begin
            tx_shift <= target_data_out;
            tx_bits_remaining <= 4'd8;
            tx_active <= 1'b1;
        end
    end
end

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        rx_shift <= '0;
        rx_bit_count <= '0;
        target_data_in <= '0;
        target_data_in_valid <= 1'b0;
    end else begin
        target_data_in_valid <= 1'b0;

        if (bus_data_in_valid && !tx_active) begin
            rx_shift[rx_bit_count] = bus_data_in;

            if (rx_bit_count == 3'd7) begin
                target_data_in <= rx_shift;
                target_data_in_valid <= 1'b1;
                rx_bit_count <= 3'd0;
                rx_shift <= '0;
            end else begin
                rx_bit_count <= rx_bit_count + 3'd1;
            end
        end
    end
end

endmodule
